module car_generator (clk,update,rst,xCount,yCount,traffic);	//this module actually generates individual lanes of traffic that move from one side of the screen to the other
input clk,rst,update;

input [9:0]xCount;
input [9:0]yCount;
wire [9:0] xCount;
wire [9:0] yCount;


output [114:0]traffic; //there are 15 lanes of traffic that each need to move at independent rates in independent directions (thus they are independent objects)
//lane 1 (top lane, 10 cars) traffic 0-9
assign traffic[0] = lane1c0;
assign traffic[1] = lane1c1;
assign traffic[2] = lane1c2;
assign traffic[3] = lane1c3;
assign traffic[4] = lane1c4;
assign traffic[5] = lane1c5;
assign traffic[6] = lane1c6;
assign traffic[7] = lane1c7;
assign traffic[8] = lane1c8;
assign traffic[9] = lane1c9;
//lane 2 (11 cars) traffic 10-20
assign traffic[10] = lane2c0;
assign traffic[11] = lane2c1;
assign traffic[12] = lane2c2;
assign traffic[13] = lane2c3;
assign traffic[14] = lane2c4;
assign traffic[15] = lane2c5;
assign traffic[16] = lane2c6;
assign traffic[17] = lane2c7;
assign traffic[18] = lane2c8;
assign traffic[19] = lane2c9;
assign traffic[20] = lane2c10;
//lane 3 (9 cars) traffic 21-29
assign traffic[21] = lane3c0;
assign traffic[22] = lane3c1;
assign traffic[23] = lane3c2;
assign traffic[24] = lane3c3;
assign traffic[25] = lane3c4;
assign traffic[26] = lane3c5;
assign traffic[27] = lane3c6;
assign traffic[28] = lane3c7;
assign traffic[29] = lane3c8;
//lane 4 (6 cars) taffic 30-35
assign traffic[30] = lane4c0;
assign traffic[31] = lane4c1;
assign traffic[32] = lane4c2;
assign traffic[33] = lane4c3;
assign traffic[34] = lane4c4;
assign traffic[35] = lane4c5;
//lane 5 (9 cars) taffic 36-45
assign traffic[36] = lane5c0;
assign traffic[37] = lane5c1;
assign traffic[38] = lane5c2;
assign traffic[39] = lane5c3;
assign traffic[40] = lane5c4;
assign traffic[41] = lane5c5;
assign traffic[42] = lane5c6;
assign traffic[43] = lane5c7;
assign traffic[44] = lane5c8;
//lane 6 (13 cars) traffic 45-57
assign traffic[45] = lane6c0;
assign traffic[46] = lane6c1;
assign traffic[47] = lane6c2;
assign traffic[48] = lane6c3;
assign traffic[49] = lane6c4;
assign traffic[50] = lane6c5;
assign traffic[51] = lane6c6;
assign traffic[52] = lane6c7;
assign traffic[53] = lane6c8;
assign traffic[54] = lane6c9;
assign traffic[55] = lane6c10;
assign traffic[56] = lane6c11;
assign traffic[57] = lane6c12;
//lane 7 (7 cars) traffic 58-64
assign traffic[58] = lane7c0;
assign traffic[59] = lane7c1;
assign traffic[60] = lane7c2;
assign traffic[61] = lane7c3;
assign traffic[62] = lane7c4;
assign traffic[63] = lane7c5;
assign traffic[64] = lane7c6;
//lane 8 (1 car) traffic 65
assign traffic[65] = lane8c0;
//lane 9 (6 cars) traffic 66-71
assign traffic[66] = lane9c0;
assign traffic[67] = lane9c1;
assign traffic[68] = lane9c2;
assign traffic[69] = lane9c3;
assign traffic[70] = lane9c4;
assign traffic[71] = lane9c5;
//lane 10 (10 cars) traffic 72-81
assign traffic[72] = lane10c0;
assign traffic[73] = lane10c1;
assign traffic[74] = lane10c2;
assign traffic[75] = lane10c3;
assign traffic[76] = lane10c4;
assign traffic[77] = lane10c5;
assign traffic[78] = lane10c6;
assign traffic[79] = lane10c7;
assign traffic[80] = lane10c8;
assign traffic[81] = lane10c9;
//lane 11 (9 cars) traffic 82-90
assign traffic[82] = lane11c0;
assign traffic[83] = lane11c1;
assign traffic[84] = lane11c2;
assign traffic[85] = lane11c3;
assign traffic[86] = lane11c4;
assign traffic[87] = lane11c5;
assign traffic[88] = lane11c6;
assign traffic[89] = lane11c7;
assign traffic[90] = lane11c8;
//lane 12 (6 cars) traffic 91-96
assign traffic[91] = lane12c0;
assign traffic[92] = lane12c1;
assign traffic[93] = lane12c2;
assign traffic[94] = lane12c3;
assign traffic[95] = lane12c4;
assign traffic[96] = lane12c5;
//lane 13 (6 cars) traffic 97-102
assign traffic[97] = lane13c0;
assign traffic[98] = lane13c1;
assign traffic[99] = lane13c2;
assign traffic[100] = lane13c3;
assign traffic[101] = lane13c4;
assign traffic[102] = lane13c5;
//lane 14 (5 cars) traffic 103-107
assign traffic[103] = lane14c0;
assign traffic[104] = lane14c1;
assign traffic[105] = lane14c2;
assign traffic[106] = lane14c3;
assign traffic[107] = lane14c4;
//lane 15 (bottom/first lane) traffic 108-115
assign traffic[108] = lane15c0;
assign traffic[109] = lane15c1;
assign traffic[110] = lane15c2;
assign traffic[111] = lane15c3;
assign traffic[112] = lane15c4;
assign traffic[113] = lane15c5;
assign traffic[114] = lane15c6;


//lane 1 
reg lane1c0;
reg lane1c1;
reg lane1c2;
reg lane1c3;
reg lane1c4;
reg lane1c5;
reg lane1c6;
reg lane1c7;
reg lane1c8;
reg lane1c9;
//lane 2 
reg lane2c0;
reg lane2c1;
reg lane2c2;
reg lane2c3;
reg lane2c4;
reg lane2c5;
reg lane2c6;
reg lane2c7;
reg lane2c8;
reg lane2c9;
reg lane2c10;
//lane 3 
reg lane3c0;
reg lane3c1;
reg lane3c2;
reg lane3c3;
reg lane3c4;
reg lane3c5;
reg lane3c6;
reg lane3c7;
reg lane3c8;
//lane 4 
reg lane4c0;
reg lane4c1;
reg lane4c2;
reg lane4c3;
reg lane4c4;
reg lane4c5;
//lane 5
reg lane5c0;
reg lane5c1;
reg lane5c2;
reg lane5c3;
reg lane5c4;
reg lane5c5;
reg lane5c6;
reg lane5c7;
reg lane5c8;
//lane 6
reg lane6c0;
reg lane6c1;
reg lane6c2;
reg lane6c3;
reg lane6c4;
reg lane6c5;
reg lane6c6;
reg lane6c7;
reg lane6c8;
reg lane6c9;
reg lane6c10;
reg lane6c11;
reg lane6c12;
//lane 7
reg lane7c0;
reg lane7c1;
reg lane7c2;
reg lane7c3;
reg lane7c4;
reg lane7c5;
reg lane7c6;
//lane 8
reg lane8c0;
//lane 9
reg lane9c0;
reg lane9c1;
reg lane9c2;
reg lane9c3;
reg lane9c4;
reg lane9c5;
//lane 10
reg lane10c0;
reg lane10c1;
reg lane10c2;
reg lane10c3;
reg lane10c4;
reg lane10c5;
reg lane10c6;
reg lane10c7;
reg lane10c8;
reg lane10c9;
//lane 11
reg lane11c0;
reg lane11c1;
reg lane11c2;
reg lane11c3;
reg lane11c4;
reg lane11c5;
reg lane11c6;
reg lane11c7;
reg lane11c8;
//lane 12
reg lane12c0;
reg lane12c1;
reg lane12c2;
reg lane12c3;
reg lane12c4;
reg lane12c5;
//lane 13
reg lane13c0;
reg lane13c1;
reg lane13c2;
reg lane13c3;
reg lane13c4;
reg lane13c5;
//lane 14
reg lane14c0;
reg lane14c1;
reg lane14c2;
reg lane14c3;
reg lane14c4;
//lane 15
reg lane15c0;
reg lane15c1;
reg lane15c2;
reg lane15c3;
reg lane15c4;
reg lane15c5;
reg lane15c6;

//lane 1 (top lane)
reg [9:0] lane1c0X [0:31];
reg [8:0] lane1c0Y [0:31];
reg [9:0] lane1c1X [0:31];
reg [8:0] lane1c1Y [0:31];
reg [9:0] lane1c2X [0:31];
reg [8:0] lane1c2Y [0:31];
reg [9:0] lane1c3X [0:31];
reg [8:0] lane1c3Y [0:31];
reg [9:0] lane1c4X [0:31];
reg [8:0] lane1c4Y [0:31];
reg [9:0] lane1c5X [0:31];
reg [8:0] lane1c5Y [0:31];
reg [9:0] lane1c6X [0:31];
reg [8:0] lane1c6Y [0:31];
reg [9:0] lane1c7X [0:31];
reg [8:0] lane1c7Y [0:31];
reg [9:0] lane1c8X [0:31];
reg [8:0] lane1c8Y [0:31];
reg [9:0] lane1c9X [0:31];
reg [8:0] lane1c9Y [0:31];
//lane 2 
reg [9:0] lane2c0X [0:31];
reg [8:0] lane2c0Y [0:31];
reg [9:0] lane2c1X [0:31];
reg [8:0] lane2c1Y [0:31];
reg [9:0] lane2c2X [0:31];
reg [8:0] lane2c2Y [0:31];
reg [9:0] lane2c3X [0:31];
reg [8:0] lane2c3Y [0:31];
reg [9:0] lane2c4X [0:31];
reg [8:0] lane2c4Y [0:31];
reg [9:0] lane2c5X [0:31];
reg [8:0] lane2c5Y [0:31];
reg [9:0] lane2c6X [0:31];
reg [8:0] lane2c6Y [0:31];
reg [9:0] lane2c7X [0:31];
reg [8:0] lane2c7Y [0:31];
reg [9:0] lane2c8X [0:31];
reg [8:0] lane2c8Y [0:31];
reg [9:0] lane2c9X [0:31];
reg [8:0] lane2c9Y [0:31];
reg [9:0] lane2c10X [0:31];
reg [8:0] lane2c10Y [0:31];
//lane 3 
reg [9:0] lane3c0X [0:31];
reg [8:0] lane3c0Y [0:31];
reg [9:0] lane3c1X [0:31];
reg [8:0] lane3c1Y [0:31];
reg [9:0] lane3c2X [0:31];
reg [8:0] lane3c2Y [0:31];
reg [9:0] lane3c3X [0:31];
reg [8:0] lane3c3Y [0:31];
reg [9:0] lane3c4X [0:31];
reg [8:0] lane3c4Y [0:31];
reg [9:0] lane3c5X [0:31];
reg [8:0] lane3c5Y [0:31];
reg [9:0] lane3c6X [0:31];
reg [8:0] lane3c6Y [0:31];
reg [9:0] lane3c7X [0:31];
reg [8:0] lane3c7Y [0:31];
reg [9:0] lane3c8X [0:31];
reg [8:0] lane3c8Y [0:31];
//lane 4 
reg [9:0] lane4c0X [0:31];
reg [8:0] lane4c0Y [0:31];
reg [9:0] lane4c1X [0:31];
reg [8:0] lane4c1Y [0:31];
reg [9:0] lane4c2X [0:31];
reg [8:0] lane4c2Y [0:31];
reg [9:0] lane4c3X [0:31];
reg [8:0] lane4c3Y [0:31];
reg [9:0] lane4c4X [0:31];
reg [8:0] lane4c4Y [0:31];
reg [9:0] lane4c5X [0:31];
reg [8:0] lane4c5Y [0:31];
//lane 5
reg [9:0] lane5c0X [0:31];
reg [8:0] lane5c0Y [0:31];
reg [9:0] lane5c1X [0:31];
reg [8:0] lane5c1Y [0:31];
reg [9:0] lane5c2X [0:31];
reg [8:0] lane5c2Y [0:31];
reg [9:0] lane5c3X [0:31];
reg [8:0] lane5c3Y [0:31];
reg [9:0] lane5c4X [0:31];
reg [8:0] lane5c4Y [0:31];
reg [9:0] lane5c5X [0:31];
reg [8:0] lane5c5Y [0:31];
reg [9:0] lane5c6X [0:31];
reg [8:0] lane5c6Y [0:31];
reg [9:0] lane5c7X [0:31];
reg [8:0] lane5c7Y [0:31];
reg [9:0] lane5c8X [0:31];
reg [8:0] lane5c8Y [0:31];
//lane 6
reg [9:0] lane6c0X [0:31];
reg [8:0] lane6c0Y [0:31];
reg [9:0] lane6c1X [0:31];
reg [8:0] lane6c1Y [0:31];
reg [9:0] lane6c2X [0:31];
reg [8:0] lane6c2Y [0:31];
reg [9:0] lane6c3X [0:31];
reg [8:0] lane6c3Y [0:31];
reg [9:0] lane6c4X [0:31];
reg [8:0] lane6c4Y [0:31];
reg [9:0] lane6c5X [0:31];
reg [8:0] lane6c5Y [0:31];
reg [9:0] lane6c6X [0:31];
reg [8:0] lane6c6Y [0:31];
reg [9:0] lane6c7X [0:31];
reg [8:0] lane6c7Y [0:31];
reg [9:0] lane6c8X [0:31];
reg [8:0] lane6c8Y [0:31];
reg [9:0] lane6c9X [0:31];
reg [8:0] lane6c9Y [0:31];
reg [9:0] lane6c10X [0:31];
reg [8:0] lane6c10Y [0:31];
reg [9:0] lane6c11X [0:31];
reg [8:0] lane6c11Y [0:31];
reg [9:0] lane6c12X [0:31];
reg [8:0] lane6c12Y [0:31];
//lane 7
reg [9:0] lane7c0X [0:31];
reg [8:0] lane7c0Y [0:31];
reg [9:0] lane7c1X [0:31];
reg [8:0] lane7c1Y [0:31];
reg [9:0] lane7c2X [0:31];
reg [8:0] lane7c2Y [0:31];
reg [9:0] lane7c3X [0:31];
reg [8:0] lane7c3Y [0:31];
reg [9:0] lane7c4X [0:31];
reg [8:0] lane7c4Y [0:31];
reg [9:0] lane7c5X [0:31];
reg [8:0] lane7c5Y [0:31];
reg [9:0] lane7c6X [0:31];
reg [8:0] lane7c6Y [0:31];
//lane 8
reg [9:0] lane8c0X [0:31];
reg [8:0] lane8c0Y [0:31];
//lane 9
reg [9:0] lane9c0X [0:31];
reg [8:0] lane9c0Y [0:31];
reg [9:0] lane9c1X [0:31];
reg [8:0] lane9c1Y [0:31];
reg [9:0] lane9c2X [0:31];
reg [8:0] lane9c2Y [0:31];
reg [9:0] lane9c3X [0:31];
reg [8:0] lane9c3Y [0:31];
reg [9:0] lane9c4X [0:31];
reg [8:0] lane9c4Y [0:31];
reg [9:0] lane9c5X [0:31];
reg [8:0] lane9c5Y [0:31];
//lane 10
reg [9:0] lane10c0X [0:31];
reg [8:0] lane10c0Y [0:31];
reg [9:0] lane10c1X [0:31];
reg [8:0] lane10c1Y [0:31];
reg [9:0] lane10c2X [0:31];
reg [8:0] lane10c2Y [0:31];
reg [9:0] lane10c3X [0:31];
reg [8:0] lane10c3Y [0:31];
reg [9:0] lane10c4X [0:31];
reg [8:0] lane10c4Y [0:31];
reg [9:0] lane10c5X [0:31];
reg [8:0] lane10c5Y [0:31];
reg [9:0] lane10c6X [0:31];
reg [8:0] lane10c6Y [0:31];
reg [9:0] lane10c7X [0:31];
reg [8:0] lane10c7Y [0:31];
reg [9:0] lane10c8X [0:31];
reg [8:0] lane10c8Y [0:31];
reg [9:0] lane10c9X [0:31];
reg [8:0] lane10c9Y [0:31];
//lane 11
reg [9:0] lane11c0X [0:31];
reg [8:0] lane11c0Y [0:31];
reg [9:0] lane11c1X [0:31];
reg [8:0] lane11c1Y [0:31];
reg [9:0] lane11c2X [0:31];
reg [8:0] lane11c2Y [0:31];
reg [9:0] lane11c3X [0:31];
reg [8:0] lane11c3Y [0:31];
reg [9:0] lane11c4X [0:31];
reg [8:0] lane11c4Y [0:31];
reg [9:0] lane11c5X [0:31];
reg [8:0] lane11c5Y [0:31];
reg [9:0] lane11c6X [0:31];
reg [8:0] lane11c6Y [0:31];
reg [9:0] lane11c7X [0:31];
reg [8:0] lane11c7Y [0:31];
reg [9:0] lane11c8X [0:31];
reg [8:0] lane11c8Y [0:31];
//lane 12
reg [9:0] lane12c0X [0:31];
reg [8:0] lane12c0Y [0:31];
reg [9:0] lane12c1X [0:31];
reg [8:0] lane12c1Y [0:31];
reg [9:0] lane12c2X [0:31];
reg [8:0] lane12c2Y [0:31];
reg [9:0] lane12c3X [0:31];
reg [8:0] lane12c3Y [0:31];
reg [9:0] lane12c4X [0:31];
reg [8:0] lane12c4Y [0:31];
reg [9:0] lane12c5X [0:31];
reg [8:0] lane12c5Y [0:31];
//lane 13
reg [9:0] lane13c0X [0:31];
reg [8:0] lane13c0Y [0:31];
reg [9:0] lane13c1X [0:31];
reg [8:0] lane13c1Y [0:31];
reg [9:0] lane13c2X [0:31];
reg [8:0] lane13c2Y [0:31];
reg [9:0] lane13c3X [0:31];
reg [8:0] lane13c3Y [0:31];
reg [9:0] lane13c4X [0:31];
reg [8:0] lane13c4Y [0:31];
reg [9:0] lane13c5X [0:31];
reg [8:0] lane13c5Y [0:31];
//lane 14
reg [9:0] lane14c0X [0:31];
reg [8:0] lane14c0Y [0:31];
reg [9:0] lane14c1X [0:31];
reg [8:0] lane14c1Y [0:31];
reg [9:0] lane14c2X [0:31];
reg [8:0] lane14c2Y [0:31];
reg [9:0] lane14c3X [0:31];
reg [8:0] lane14c3Y [0:31];
reg [9:0] lane14c4X [0:31];
reg [8:0] lane14c4Y [0:31];
//lane 15
reg [9:0] lane15c0X [0:31];
reg [8:0] lane15c0Y [0:31];
reg [9:0] lane15c1X [0:31];
reg [8:0] lane15c1Y [0:31];
reg [9:0] lane15c2X [0:31];
reg [8:0] lane15c2Y [0:31];
reg [9:0] lane15c3X [0:31];
reg [8:0] lane15c3Y [0:31];
reg [9:0] lane15c4X [0:31];
reg [8:0] lane15c4Y [0:31];
reg [9:0] lane15c5X [0:31];
reg [8:0] lane15c5Y [0:31];
reg [9:0] lane15c6X [0:31];
reg [8:0] lane15c6Y [0:31];


//controls the size of the "cars"
always@(posedge clk) 
	begin	
		//lane 1 (top lane, 10 cars)
		lane1c0 <= (xCount > lane1c0X[0] && xCount < (lane1c0X[0]+17)) && (yCount > lane1c0Y[0] && yCount < (lane1c0Y[0]+17));
		lane1c1 <= (xCount > lane1c1X[0] && xCount < (lane1c1X[0]+30)) && (yCount > lane1c1Y[0] && yCount < (lane1c1Y[0]+17));
		lane1c2 <= (xCount > lane1c2X[0] && xCount < (lane1c2X[0]+17)) && (yCount > lane1c2Y[0] && yCount < (lane1c2Y[0]+17));
		lane1c3 <= (xCount > lane1c3X[0] && xCount < (lane1c3X[0]+25)) && (yCount > lane1c3Y[0] && yCount < (lane1c3Y[0]+17));
		lane1c4 <= (xCount > lane1c4X[0] && xCount < (lane1c4X[0]+17)) && (yCount > lane1c4Y[0] && yCount < (lane1c4Y[0]+17));
		lane1c5 <= (xCount > lane1c5X[0] && xCount < (lane1c5X[0]+27)) && (yCount > lane1c5Y[0] && yCount < (lane1c5Y[0]+17));
		lane1c6 <= (xCount > lane1c6X[0] && xCount < (lane1c6X[0]+17)) && (yCount > lane1c6Y[0] && yCount < (lane1c6Y[0]+17));
		lane1c7 <= (xCount > lane1c7X[0] && xCount < (lane1c7X[0]+33)) && (yCount > lane1c7Y[0] && yCount < (lane1c7Y[0]+17));
		lane1c8 <= (xCount > lane1c8X[0] && xCount < (lane1c8X[0]+17)) && (yCount > lane1c8Y[0] && yCount < (lane1c8Y[0]+17));
		lane1c9 <= (xCount > lane1c9X[0] && xCount < (lane1c9X[0]+31)) && (yCount > lane1c9Y[0] && yCount < (lane1c9Y[0]+17));
		
		//lane 2 (11 cars)
		lane2c0 <= (xCount > lane2c0X[0] && xCount < (lane2c0X[0]+17)) && (yCount > lane2c0Y[0] && yCount < (lane2c0Y[0]+17));
		lane2c1 <= (xCount > lane2c1X[0] && xCount < (lane2c1X[0]+17)) && (yCount > lane2c1Y[0] && yCount < (lane2c1Y[0]+17));
		lane2c2 <= (xCount > lane2c2X[0] && xCount < (lane2c2X[0]+26)) && (yCount > lane2c2Y[0] && yCount < (lane2c2Y[0]+17));
		lane2c3 <= (xCount > lane2c3X[0] && xCount < (lane2c3X[0]+17)) && (yCount > lane2c3Y[0] && yCount < (lane2c3Y[0]+17));
		lane2c4 <= (xCount > lane2c4X[0] && xCount < (lane2c4X[0]+17)) && (yCount > lane2c4Y[0] && yCount < (lane2c4Y[0]+17));
		lane2c5 <= (xCount > lane2c5X[0] && xCount < (lane2c5X[0]+17)) && (yCount > lane2c5Y[0] && yCount < (lane2c5Y[0]+17));
		lane2c6 <= (xCount > lane2c6X[0] && xCount < (lane2c6X[0]+17)) && (yCount > lane2c6Y[0] && yCount < (lane2c6Y[0]+17));
		lane2c7 <= (xCount > lane2c7X[0] && xCount < (lane2c7X[0]+17)) && (yCount > lane2c7Y[0] && yCount < (lane2c7Y[0]+17));
		lane2c8 <= (xCount > lane2c8X[0] && xCount < (lane2c8X[0]+17)) && (yCount > lane2c8Y[0] && yCount < (lane2c8Y[0]+17));
		lane2c9 <= (xCount > lane2c9X[0] && xCount < (lane2c9X[0]+17)) && (yCount > lane2c9Y[0] && yCount < (lane2c9Y[0]+17));
		lane2c10 <= (xCount > lane2c10X[0] && xCount < (lane2c10X[0]+17)) && (yCount > lane2c10Y[0] && yCount < (lane2c10Y[0]+17));

		//lane 3 (9 cars)
		lane3c0 <= (xCount > lane3c0X[0] && xCount < (lane3c0X[0]+17)) && (yCount > lane3c0Y[0] && yCount < (lane3c0Y[0]+17));
		lane3c1 <= (xCount > lane3c1X[0] && xCount < (lane3c1X[0]+17)) && (yCount > lane3c1Y[0] && yCount < (lane3c1Y[0]+17));
		lane3c2 <= (xCount > lane3c2X[0] && xCount < (lane3c2X[0]+17)) && (yCount > lane3c2Y[0] && yCount < (lane3c2Y[0]+17));
		lane3c3 <= (xCount > lane3c3X[0] && xCount < (lane3c3X[0]+17)) && (yCount > lane3c3Y[0] && yCount < (lane3c3Y[0]+17));
		lane3c4 <= (xCount > lane3c4X[0] && xCount < (lane3c4X[0]+17)) && (yCount > lane3c4Y[0] && yCount < (lane3c4Y[0]+17));
		lane3c5 <= (xCount > lane3c5X[0] && xCount < (lane3c5X[0]+17)) && (yCount > lane3c5Y[0] && yCount < (lane3c5Y[0]+17));
		lane3c6 <= (xCount > lane3c6X[0] && xCount < (lane3c6X[0]+17)) && (yCount > lane3c6Y[0] && yCount < (lane3c6Y[0]+17));
		lane3c7 <= (xCount > lane3c7X[0] && xCount < (lane3c7X[0]+17)) && (yCount > lane3c7Y[0] && yCount < (lane3c7Y[0]+17));
		lane3c8 <= (xCount > lane3c8X[0] && xCount < (lane3c8X[0]+17)) && (yCount > lane3c8Y[0] && yCount < (lane3c8Y[0]+17));
		
		//lane 4 (6 cars)
		lane4c0 <= (xCount > lane4c0X[0] && xCount < (lane4c0X[0]+17)) && (yCount > lane4c0Y[0] && yCount < (lane4c0Y[0]+17));
		lane4c1 <= (xCount > lane4c1X[0] && xCount < (lane4c1X[0]+40)) && (yCount > lane4c1Y[0] && yCount < (lane4c1Y[0]+17));
		lane4c2 <= (xCount > lane4c2X[0] && xCount < (lane4c2X[0]+35)) && (yCount > lane4c2Y[0] && yCount < (lane4c2Y[0]+17));
		lane4c3 <= (xCount > lane4c3X[0] && xCount < (lane4c3X[0]+25)) && (yCount > lane4c3Y[0] && yCount < (lane4c3Y[0]+17));
		lane4c4 <= (xCount > lane4c4X[0] && xCount < (lane4c4X[0]+17)) && (yCount > lane4c4Y[0] && yCount < (lane4c4Y[0]+17));
		lane4c5 <= (xCount > lane4c5X[0] && xCount < (lane4c5X[0]+30)) && (yCount > lane4c5Y[0] && yCount < (lane4c5Y[0]+17));
		
		//lane 5
		lane5c0 <= (xCount > lane5c0X[0] && xCount < (lane5c0X[0]+17)) && (yCount > lane5c0Y[0] && yCount < (lane5c0Y[0]+17));
		lane5c1 <= (xCount > lane5c1X[0] && xCount < (lane5c1X[0]+17)) && (yCount > lane5c1Y[0] && yCount < (lane5c1Y[0]+17));
		lane5c2 <= (xCount > lane5c2X[0] && xCount < (lane5c2X[0]+17)) && (yCount > lane5c2Y[0] && yCount < (lane5c2Y[0]+17));
		lane5c3 <= (xCount > lane5c3X[0] && xCount < (lane5c3X[0]+17)) && (yCount > lane5c3Y[0] && yCount < (lane5c3Y[0]+17));
		lane5c4 <= (xCount > lane5c4X[0] && xCount < (lane5c4X[0]+17)) && (yCount > lane5c4Y[0] && yCount < (lane5c4Y[0]+17));
		lane5c5 <= (xCount > lane5c5X[0] && xCount < (lane5c5X[0]+17)) && (yCount > lane5c5Y[0] && yCount < (lane5c5Y[0]+17));
		lane5c6 <= (xCount > lane5c6X[0] && xCount < (lane5c6X[0]+17)) && (yCount > lane5c6Y[0] && yCount < (lane5c6Y[0]+17));
		lane5c7 <= (xCount > lane5c7X[0] && xCount < (lane5c7X[0]+17)) && (yCount > lane5c7Y[0] && yCount < (lane5c7Y[0]+17));
		lane5c8 <= (xCount > lane5c8X[0] && xCount < (lane5c8X[0]+17)) && (yCount > lane5c8Y[0] && yCount < (lane5c8Y[0]+17));
		
		//lane 6
		lane6c0 <= (xCount > lane6c0X[0] && xCount < (lane6c0X[0]+17)) && (yCount > lane6c0Y[0] && yCount < (lane6c0Y[0]+17));
		lane6c1 <= (xCount > lane6c1X[0] && xCount < (lane6c1X[0]+17)) && (yCount > lane6c1Y[0] && yCount < (lane6c1Y[0]+17));
		lane6c2 <= (xCount > lane6c2X[0] && xCount < (lane6c2X[0]+17)) && (yCount > lane6c2Y[0] && yCount < (lane6c2Y[0]+17));
		lane6c3 <= (xCount > lane6c3X[0] && xCount < (lane6c3X[0]+17)) && (yCount > lane6c3Y[0] && yCount < (lane6c3Y[0]+17));
		lane6c4 <= (xCount > lane6c4X[0] && xCount < (lane6c4X[0]+17)) && (yCount > lane6c4Y[0] && yCount < (lane6c4Y[0]+17));
		lane6c5 <= (xCount > lane6c5X[0] && xCount < (lane6c5X[0]+17)) && (yCount > lane6c5Y[0] && yCount < (lane6c5Y[0]+17));
		lane6c6 <= (xCount > lane6c6X[0] && xCount < (lane6c6X[0]+17)) && (yCount > lane6c6Y[0] && yCount < (lane6c6Y[0]+17));
		lane6c7 <= (xCount > lane6c7X[0] && xCount < (lane6c7X[0]+17)) && (yCount > lane6c7Y[0] && yCount < (lane6c7Y[0]+17));
		lane6c8 <= (xCount > lane6c8X[0] && xCount < (lane6c8X[0]+17)) && (yCount > lane6c8Y[0] && yCount < (lane6c8Y[0]+17));
		lane6c9 <= (xCount > lane6c9X[0] && xCount < (lane6c9X[0]+17)) && (yCount > lane6c9Y[0] && yCount < (lane6c9Y[0]+17));
		lane6c10 <= (xCount > lane6c10X[0] && xCount < (lane6c10X[0]+17)) && (yCount > lane6c10Y[0] && yCount < (lane6c10Y[0]+17));
		lane6c11 <= (xCount > lane6c11X[0] && xCount < (lane6c11X[0]+17)) && (yCount > lane6c11Y[0] && yCount < (lane6c11Y[0]+17));
		lane6c12 <= (xCount > lane6c12X[0] && xCount < (lane6c12X[0]+17)) && (yCount > lane6c12Y[0] && yCount < (lane6c12Y[0]+17));
		
		//lane 7
		lane7c0 <= (xCount > lane7c0X[0] && xCount < (lane7c0X[0]+25)) && (yCount > lane7c0Y[0] && yCount < (lane7c0Y[0]+17));
		lane7c1 <= (xCount > lane7c1X[0] && xCount < (lane7c1X[0]+25)) && (yCount > lane7c1Y[0] && yCount < (lane7c1Y[0]+17));
		lane7c2 <= (xCount > lane7c2X[0] && xCount < (lane7c2X[0]+25)) && (yCount > lane7c2Y[0] && yCount < (lane7c2Y[0]+17));
		lane7c3 <= (xCount > lane7c3X[0] && xCount < (lane7c3X[0]+25)) && (yCount > lane7c3Y[0] && yCount < (lane7c3Y[0]+17));
		lane7c4 <= (xCount > lane7c4X[0] && xCount < (lane7c4X[0]+25)) && (yCount > lane7c4Y[0] && yCount < (lane7c4Y[0]+17));
		lane7c5 <= (xCount > lane7c5X[0] && xCount < (lane7c5X[0]+25)) && (yCount > lane7c5Y[0] && yCount < (lane7c5Y[0]+17));
		lane7c6 <= (xCount > lane7c6X[0] && xCount < (lane7c6X[0]+25)) && (yCount > lane7c6Y[0] && yCount < (lane7c6Y[0]+17));
		
		//lane 8
		lane8c0 <= (xCount > lane8c0X[0] && xCount < (lane8c0X[0]+17)) && (yCount > lane8c0Y[0] && yCount < (lane8c0Y[0]+17));
		
		//lane 9
		lane9c0 <= (xCount > lane9c0X[0] && xCount < (lane9c0X[0]+20)) && (yCount > lane9c0Y[0] && yCount < (lane9c0Y[0]+17));
		lane9c1 <= (xCount > lane9c1X[0] && xCount < (lane9c1X[0]+20)) && (yCount > lane9c1Y[0] && yCount < (lane9c1Y[0]+17));
		lane9c2 <= (xCount > lane9c2X[0] && xCount < (lane9c2X[0]+20)) && (yCount > lane9c2Y[0] && yCount < (lane9c2Y[0]+17));
		lane9c3 <= (xCount > lane9c3X[0] && xCount < (lane9c3X[0]+20)) && (yCount > lane9c3Y[0] && yCount < (lane9c3Y[0]+17));
		lane9c4 <= (xCount > lane9c4X[0] && xCount < (lane9c4X[0]+20)) && (yCount > lane9c4Y[0] && yCount < (lane9c4Y[0]+17));
		lane9c5 <= (xCount > lane9c5X[0] && xCount < (lane9c5X[0]+20)) && (yCount > lane9c5Y[0] && yCount < (lane9c5Y[0]+17));
		
		//lane 10
		lane10c0 <= (xCount > lane10c0X[0] && xCount < (lane10c0X[0]+17)) && (yCount > lane10c0Y[0] && yCount < (lane10c0Y[0]+17));
		lane10c1 <= (xCount > lane10c1X[0] && xCount < (lane10c1X[0]+17)) && (yCount > lane10c1Y[0] && yCount < (lane10c1Y[0]+17));
		lane10c2 <= (xCount > lane10c2X[0] && xCount < (lane10c2X[0]+17)) && (yCount > lane10c2Y[0] && yCount < (lane10c2Y[0]+17));
		lane10c3 <= (xCount > lane10c3X[0] && xCount < (lane10c3X[0]+17)) && (yCount > lane10c3Y[0] && yCount < (lane10c3Y[0]+17));
		lane10c4 <= (xCount > lane10c4X[0] && xCount < (lane10c4X[0]+17)) && (yCount > lane10c4Y[0] && yCount < (lane10c4Y[0]+17));
		lane10c5 <= (xCount > lane10c5X[0] && xCount < (lane10c5X[0]+17)) && (yCount > lane10c5Y[0] && yCount < (lane10c5Y[0]+17));
		lane10c6 <= (xCount > lane10c6X[0] && xCount < (lane10c6X[0]+17)) && (yCount > lane10c6Y[0] && yCount < (lane10c6Y[0]+17));
		lane10c7 <= (xCount > lane10c7X[0] && xCount < (lane10c7X[0]+17)) && (yCount > lane10c7Y[0] && yCount < (lane10c7Y[0]+17));
		lane10c8 <= (xCount > lane10c8X[0] && xCount < (lane10c8X[0]+17)) && (yCount > lane10c8Y[0] && yCount < (lane10c8Y[0]+17));
		lane10c9 <= (xCount > lane10c9X[0] && xCount < (lane10c9X[0]+17)) && (yCount > lane10c9Y[0] && yCount < (lane10c9Y[0]+17));
		
		//lane 11
		lane11c0 <= (xCount > lane11c0X[0] && xCount < (lane11c0X[0]+17)) && (yCount > lane11c0Y[0] && yCount < (lane11c0Y[0]+17));
		lane11c1 <= (xCount > lane11c1X[0] && xCount < (lane11c1X[0]+17)) && (yCount > lane11c1Y[0] && yCount < (lane11c1Y[0]+17));
		lane11c2 <= (xCount > lane11c2X[0] && xCount < (lane11c2X[0]+17)) && (yCount > lane11c2Y[0] && yCount < (lane11c2Y[0]+17));
		lane11c3 <= (xCount > lane11c3X[0] && xCount < (lane11c3X[0]+17)) && (yCount > lane11c3Y[0] && yCount < (lane11c3Y[0]+17));
		lane11c4 <= (xCount > lane11c4X[0] && xCount < (lane11c4X[0]+17)) && (yCount > lane11c4Y[0] && yCount < (lane11c4Y[0]+17));
		lane11c5 <= (xCount > lane11c5X[0] && xCount < (lane11c5X[0]+17)) && (yCount > lane11c5Y[0] && yCount < (lane11c5Y[0]+17));
		lane11c6 <= (xCount > lane11c6X[0] && xCount < (lane11c6X[0]+17)) && (yCount > lane11c6Y[0] && yCount < (lane11c6Y[0]+17));
		lane11c7 <= (xCount > lane11c7X[0] && xCount < (lane11c7X[0]+17)) && (yCount > lane11c7Y[0] && yCount < (lane11c7Y[0]+17));
		lane11c8 <= (xCount > lane11c8X[0] && xCount < (lane11c8X[0]+17)) && (yCount > lane11c8Y[0] && yCount < (lane11c8Y[0]+17));
		
		//lane 12
		lane12c0 <= (xCount > lane12c0X[0] && xCount < (lane12c0X[0]+17)) && (yCount > lane12c0Y[0] && yCount < (lane12c0Y[0]+17));
		lane12c1 <= (xCount > lane12c1X[0] && xCount < (lane12c1X[0]+17)) && (yCount > lane12c1Y[0] && yCount < (lane12c1Y[0]+17));
		lane12c2 <= (xCount > lane12c2X[0] && xCount < (lane12c2X[0]+17)) && (yCount > lane12c2Y[0] && yCount < (lane12c2Y[0]+17));
		lane12c3 <= (xCount > lane12c3X[0] && xCount < (lane12c3X[0]+17)) && (yCount > lane12c3Y[0] && yCount < (lane12c3Y[0]+17));
		lane12c4 <= (xCount > lane12c4X[0] && xCount < (lane12c4X[0]+17)) && (yCount > lane12c4Y[0] && yCount < (lane12c4Y[0]+17));
		lane12c5 <= (xCount > lane12c5X[0] && xCount < (lane12c5X[0]+17)) && (yCount > lane12c5Y[0] && yCount < (lane12c5Y[0]+17));
		
		//lane 13
		lane13c0 <= (xCount > lane13c0X[0] && xCount < (lane13c0X[0]+22)) && (yCount > lane13c0Y[0] && yCount < (lane13c0Y[0]+17));
		lane13c1 <= (xCount > lane13c1X[0] && xCount < (lane13c1X[0]+22)) && (yCount > lane13c1Y[0] && yCount < (lane13c1Y[0]+17));
		lane13c2 <= (xCount > lane13c2X[0] && xCount < (lane13c2X[0]+22)) && (yCount > lane13c2Y[0] && yCount < (lane13c2Y[0]+17));
		lane13c3 <= (xCount > lane13c3X[0] && xCount < (lane13c3X[0]+22)) && (yCount > lane13c3Y[0] && yCount < (lane13c3Y[0]+17));
		lane13c4 <= (xCount > lane13c4X[0] && xCount < (lane13c4X[0]+22)) && (yCount > lane13c4Y[0] && yCount < (lane13c4Y[0]+17));
		lane13c5 <= (xCount > lane13c5X[0] && xCount < (lane13c5X[0]+22)) && (yCount > lane13c5Y[0] && yCount < (lane13c5Y[0]+17));
		
		//lane 14
		lane14c0 <= (xCount > lane14c0X[0] && xCount < (lane14c0X[0]+30)) && (yCount > lane14c0Y[0] && yCount < (lane14c0Y[0]+17));
		lane14c1 <= (xCount > lane14c1X[0] && xCount < (lane14c1X[0]+30)) && (yCount > lane14c1Y[0] && yCount < (lane14c1Y[0]+17));
		lane14c2 <= (xCount > lane14c2X[0] && xCount < (lane14c2X[0]+30)) && (yCount > lane14c2Y[0] && yCount < (lane14c2Y[0]+17));
		lane14c3 <= (xCount > lane14c3X[0] && xCount < (lane14c3X[0]+30)) && (yCount > lane14c3Y[0] && yCount < (lane14c3Y[0]+17));
		lane14c4 <= (xCount > lane14c4X[0] && xCount < (lane14c4X[0]+30)) && (yCount > lane14c4Y[0] && yCount < (lane14c4Y[0]+17));
		
		//lane 15
		lane15c0 <= (xCount > lane15c0X[0] && xCount < (lane15c0X[0]+17)) && (yCount > lane15c0Y[0] && yCount < (lane15c0Y[0]+17));
		lane15c1 <= (xCount > lane15c1X[0] && xCount < (lane15c1X[0]+17)) && (yCount > lane15c1Y[0] && yCount < (lane15c1Y[0]+17));
		lane15c2 <= (xCount > lane15c2X[0] && xCount < (lane15c2X[0]+17)) && (yCount > lane15c2Y[0] && yCount < (lane15c2Y[0]+17));
		lane15c3 <= (xCount > lane15c3X[0] && xCount < (lane15c3X[0]+17)) && (yCount > lane15c3Y[0] && yCount < (lane15c3Y[0]+17));
		lane15c4 <= (xCount > lane15c4X[0] && xCount < (lane15c4X[0]+17)) && (yCount > lane15c4Y[0] && yCount < (lane15c4Y[0]+17));
		lane15c5 <= (xCount > lane15c5X[0] && xCount < (lane15c5X[0]+17)) && (yCount > lane15c5Y[0] && yCount < (lane15c5Y[0]+17));
		lane15c6 <= (xCount > lane15c6X[0] && xCount < (lane15c6X[0]+17)) && (yCount > lane15c6Y[0] && yCount < (lane15c6Y[0]+17));
				
	end
//	

/////lane1 control /////
always @(posedge update)
	begin
		if (rst == 1'b1)
			begin //starting position of lane1 cars				
				lane1c0X[0] <= 20;
				lane1c0Y[0] <= 74;
				lane1c1X[0] <= 90;
				lane1c1Y[0] <= 74;
				lane1c2X[0] <= 160;
				lane1c2Y[0] <= 74;
				lane1c3X[0] <= 230;
				lane1c3Y[0] <= 74;
				lane1c4X[0] <= 300;
				lane1c4Y[0] <= 74;
				lane1c5X[0] <= 370;
				lane1c5Y[0] <= 74;
				lane1c6X[0] <= 440;
				lane1c6Y[0] <= 74;
				lane1c7X[0] <= 510;
				lane1c7Y[0] <= 74;
				lane1c8X[0] <= 580;
				lane1c8Y[0] <= 74;
				lane1c9X[0] <= 610;
				lane1c9Y[0] <= 74;
			end
			
		//recycling cars back to the start of the lane
		else if (lane1c0X[0] >= 640)
			lane1c0X[0] <= 0;
		else if (lane1c1X[0] >= 640)
			lane1c1X[0] <= 0;
		else if (lane1c2X[0] >= 640)
			lane1c2X[0] <= 0;
		else if (lane1c3X[0] >= 640)
			lane1c3X[0] <= 0;
		else if (lane1c4X[0] >= 640)
			lane1c4X[0] <= 0;
		else if (lane1c5X[0] >= 640)
			lane1c5X[0] <= 0;
		else if (lane1c6X[0] >= 640)
			lane1c6X[0] <= 0;
		else if (lane1c7X[0] >= 640)
			lane1c7X[0] <= 0;
		else if (lane1c8X[0] >= 640)
			lane1c8X[0] <= 0;
		else if (lane1c9X[0] >= 640)
			lane1c9X[0] <= 0;
	
		else
			begin //rate and direction of cars
				lane1c0X[0] <= lane1c0X[0] + 2;
				lane1c1X[0] <= lane1c1X[0] + 2;
				lane1c2X[0] <= lane1c2X[0] + 2;
				lane1c3X[0] <= lane1c3X[0] + 2;
				lane1c4X[0] <= lane1c4X[0] + 2;
				lane1c5X[0] <= lane1c5X[0] + 2;
				lane1c6X[0] <= lane1c6X[0] + 2;
				lane1c7X[0] <= lane1c7X[0] + 2;
				lane1c8X[0] <= lane1c8X[0] + 2;
				lane1c9X[0] <= lane1c9X[0] + 2;	
			end
	end
//

///// lane2 control /////
always @(posedge update)
	begin
		if (rst == 1'b1) //starting positions of lane2 cars
			begin
				lane2c0X[0] <= 20;
				lane2c0Y[0] <= 99;
				lane2c1X[0] <= 90;
				lane2c1Y[0] <= 99;
				lane2c2X[0] <= 160;
				lane2c2Y[0] <= 99;
				lane2c3X[0] <= 230;
				lane2c3Y[0] <= 99;
				lane2c4X[0] <= 300;
				lane2c4Y[0] <= 99;
				lane2c5X[0] <= 370;
				lane2c5Y[0] <= 99;
				lane2c6X[0] <= 440;
				lane2c6Y[0] <= 99;
				lane2c7X[0] <= 510;
				lane2c7Y[0] <= 99;
				lane2c8X[0] <= 580;
				lane2c8Y[0] <= 99;
				lane2c9X[0] <= 610;
				lane2c9Y[0] <= 99;
				lane2c10X[0] <= 470;
				lane2c10Y[0] <= 99;
			end
			
		//recycle cars back to start of the lane
		else if (lane2c0X[0] >= 640)
			lane2c0X[0] <= 0;
		else if (lane2c1X[0] >= 640)
			lane2c1X[0] <= 0;
		else if (lane2c2X[0] >= 640)
			lane2c2X[0] <= 0;
		else if (lane2c3X[0] >= 640)
			lane2c3X[0] <= 0;
		else if (lane2c4X[0] >= 640)
			lane2c4X[0] <= 0;
		else if (lane2c5X[0] >= 640)
			lane2c5X[0] <= 0;
		else if (lane2c6X[0] >= 640)
			lane2c6X[0] <= 0;
		else if (lane2c7X[0] >= 640)
			lane2c7X[0] <= 0;
		else if (lane2c8X[0] >= 640)
			lane2c8X[0] <= 0;
		else if (lane2c9X[0] >= 640)
			lane2c9X[0] <= 0;
		else if (lane2c10X[0] >= 640)
			lane2c10X[0] <= 0;
			
		else //rate and direction of cars
			begin
				lane2c0X[0] <= lane2c0X[0] + 1;
				lane2c1X[0] <= lane2c1X[0] + 1;
				lane2c2X[0] <= lane2c2X[0] + 1;
				lane2c3X[0] <= lane2c3X[0] + 1;
				lane2c4X[0] <= lane2c4X[0] + 1;
				lane2c5X[0] <= lane2c5X[0] + 1;
				lane2c6X[0] <= lane2c6X[0] + 1;
				lane2c7X[0] <= lane2c7X[0] + 1;
				lane2c8X[0] <= lane2c8X[0] + 1;
				lane2c9X[0] <= lane2c9X[0] + 1;
				lane2c10X[0] <= lane2c10X[0] + 1;
			end
		end
//

/////lane3 control /////
always @(posedge update)
	begin
		if (rst == 1'b1)
			begin //starting position of lane3 cars
				lane3c0X[0] <= 30;
				lane3c0Y[0] <= 124;
				lane3c1X[0] <= 100;
				lane3c1Y[0] <= 124;
				lane3c2X[0] <= 170;
				lane3c2Y[0] <= 124;
				lane3c3X[0] <= 240;
				lane3c3Y[0] <= 124;
				lane3c4X[0] <= 310;
				lane3c4Y[0] <= 124;
				lane3c5X[0] <= 380;
				lane3c5Y[0] <= 124;
				lane3c6X[0] <= 450;
				lane3c6Y[0] <= 124;
				lane3c7X[0] <= 520;
				lane3c7Y[0] <= 124;
				lane3c8X[0] <= 580;
				lane3c8Y[0] <= 124;
			end
		//recycling cars back to the start of the lane
		else if (lane3c0X[0] == 0)
			lane3c0X[0] <= 640;
		else if (lane3c1X[0] == 0)
			lane3c1X[0] <= 640;
		else if (lane3c2X[0] == 0)
			lane3c2X[0] <= 640;
		else if (lane3c3X[0] == 0)
			lane3c3X[0] <= 640;
		else if (lane3c4X[0] == 0)
			lane3c4X[0] <= 640;
		else if (lane3c5X[0] == 0)
			lane3c5X[0] <= 640;
		else if (lane3c6X[0] == 0)
			lane3c6X[0] <= 640;
		else if (lane3c7X[0] == 0)
			lane3c7X[0] <= 640;
		else if (lane3c8X[0] == 0)
			lane3c8X[0] <= 640;
		else
			begin //rate and direction of cars
				lane3c0X[0] <= lane3c0X[0] - 1;
				lane3c1X[0] <= lane3c1X[0] - 1;
				lane3c2X[0] <= lane3c2X[0] - 1;
				lane3c3X[0] <= lane3c3X[0] - 1;
				lane3c4X[0] <= lane3c4X[0] - 1;
				lane3c5X[0] <= lane3c5X[0] - 1;
				lane3c6X[0] <= lane3c6X[0] - 1;
				lane3c7X[0] <= lane3c7X[0] - 1;
				lane3c8X[0] <= lane3c8X[0] - 1;
			end
	end
//

/////lane4 control /////
always @(posedge update)
	begin
		if (rst == 1'b1)
			begin //starting position of lane4 cars				
				lane4c0X[0] <= 20;
				lane4c0Y[0] <= 149;
				lane4c1X[0] <= 90;
				lane4c1Y[0] <= 149;
				lane4c2X[0] <= 210;
				lane4c2Y[0] <= 149;
				lane4c3X[0] <= 330;
				lane4c3Y[0] <= 149;
				lane4c4X[0] <= 450;
				lane4c4Y[0] <= 149;
				lane4c5X[0] <= 570;
				lane4c5Y[0] <= 149;
				
			end
			
		//recycling cars back to the start of the lane
		else if (lane4c0X[0] >= 640)
			lane4c0X[0] <= 0;
		else if (lane4c1X[0] >= 640)
			lane4c1X[0] <= 0;
		else if (lane4c2X[0] >= 640)
			lane4c2X[0] <= 0;
		else if (lane4c3X[0] >= 640)
			lane4c3X[0] <= 0;
		else if (lane4c4X[0] >= 640)
			lane4c4X[0] <= 0;
		else if (lane4c5X[0] >= 640)
			lane4c5X[0] <= 0;
			
		else
			begin //rate and direction of cars
				lane4c0X[0] <= lane4c0X[0] + 3;
				lane4c1X[0] <= lane4c1X[0] + 3;
				lane4c2X[0] <= lane4c2X[0] + 3;
				lane4c3X[0] <= lane4c3X[0] + 3;
				lane4c4X[0] <= lane4c4X[0] + 3;
				lane4c5X[0] <= lane4c5X[0] + 3;
					
			end
	end
//

/////lane5 control /////
always @(posedge update)
	begin
		if (rst == 1'b1)
			begin //starting position of lane5 cars
				lane5c0X[0] <= 20;
				lane5c0Y[0] <= 174;
				lane5c1X[0] <= 90;
				lane5c1Y[0] <= 174;
				lane5c2X[0] <= 160;
				lane5c2Y[0] <= 174;
				lane5c3X[0] <= 230;
				lane5c3Y[0] <= 174;
				lane5c4X[0] <= 300;
				lane5c4Y[0] <= 174;
				lane5c5X[0] <= 370;
				lane5c5Y[0] <= 174;
				lane5c6X[0] <= 440;
				lane5c6Y[0] <= 174;
				lane5c7X[0] <= 510;
				lane5c7Y[0] <= 174;
				lane5c8X[0] <= 580;
				lane5c8Y[0] <= 174;
			end
		//recycling cars back to the start of the lane
		else if (lane5c0X[0] == 0)
			lane5c0X[0] <= 640;
		else if (lane5c1X[0] == 0)
			lane5c1X[0] <= 640;
		else if (lane5c2X[0] == 0)
			lane5c2X[0] <= 640;
		else if (lane5c3X[0] == 0)
			lane5c3X[0] <= 640;
		else if (lane5c4X[0] == 0)
			lane5c4X[0] <= 640;
		else if (lane5c5X[0] == 0)
			lane5c5X[0] <= 640;
		else if (lane5c6X[0] == 0)
			lane5c6X[0] <= 640;
		else if (lane5c7X[0] == 0)
			lane5c7X[0] <= 640;
		else if (lane5c8X[0] == 0)
			lane5c8X[0] <= 640;
		else
			begin //rate and direction of cars
				lane5c0X[0] <= lane5c0X[0] - 2;
				lane5c1X[0] <= lane5c1X[0] - 2;
				lane5c2X[0] <= lane5c2X[0] - 2;
				lane5c3X[0] <= lane5c3X[0] - 2;
				lane5c4X[0] <= lane5c4X[0] - 2;
				lane5c5X[0] <= lane5c5X[0] - 2;
				lane5c6X[0] <= lane5c6X[0] - 2;
				lane5c7X[0] <= lane5c7X[0] - 2;
				lane5c8X[0] <= lane5c8X[0] - 2;
			end
	end
//

/////lane6 control /////
always @(posedge update)
	begin
		if (rst == 1'b1)
			begin //starting position of lane6 cars
				lane6c0X[0] <= 20;
				lane6c0Y[0] <= 199;
				lane6c1X[0] <= 90;
				lane6c1Y[0] <= 199;
				lane6c2X[0] <= 160;
				lane6c2Y[0] <= 199;
				lane6c3X[0] <= 230;
				lane6c3Y[0] <= 199;
				lane6c4X[0] <= 300;
				lane6c4Y[0] <= 199;
				lane6c5X[0] <= 370;
				lane6c5Y[0] <= 199;
				lane6c6X[0] <= 440;
				lane6c6Y[0] <= 199;
				lane6c7X[0] <= 510;
				lane6c7Y[0] <= 199;
				lane6c8X[0] <= 580;
				lane6c8Y[0] <= 199;
				lane6c9X[0] <= 610;
				lane6c9Y[0] <= 199;
				lane6c10X[0] <= 470;
				lane6c10Y[0] <= 199;
				lane6c11X[0] <= 260;
				lane6c11Y[0] <= 199;
				lane6c12X[0] <= 130;
				lane6c12Y[0] <= 199;
				
			end
		//recycling cars back to the start of the lane
		else if (lane6c0X[0] == 0)
			lane6c0X[0] <= 640;
		else if (lane6c1X[0] == 0)
			lane6c1X[0] <= 640;
		else if (lane6c2X[0] == 0)
			lane6c2X[0] <= 640;
		else if (lane6c3X[0] == 0)
			lane6c3X[0] <= 640;
		else if (lane6c4X[0] == 0)
			lane6c4X[0] <= 640;
		else if (lane6c5X[0] == 0)
			lane6c5X[0] <= 640;
		else if (lane6c6X[0] == 0)
			lane6c6X[0] <= 640;
		else if (lane6c7X[0] == 0)
			lane6c7X[0] <= 640;
		else if (lane6c8X[0] == 0)
			lane6c8X[0] <= 640;
		else if (lane6c9X[0] == 0)
			lane6c9X[0] <= 640;
		else if (lane6c10X[0] == 0)
			lane6c10X[0] <= 640;
		else if (lane6c11X[0] == 0)
			lane6c11X[0] <= 640;
		else if (lane6c12X[0] == 0)
			lane6c12X[0] <= 640;
	
		else
			begin //rate and direction of cars
				lane6c0X[0] <= lane6c0X[0] - 1;
				lane6c1X[0] <= lane6c1X[0] - 1;
				lane6c2X[0] <= lane6c2X[0] - 1;
				lane6c3X[0] <= lane6c3X[0] - 1;
				lane6c4X[0] <= lane6c4X[0] - 1;
				lane6c5X[0] <= lane6c5X[0] - 1;
				lane6c6X[0] <= lane6c6X[0] - 1;
				lane6c7X[0] <= lane6c7X[0] - 1;
				lane6c8X[0] <= lane6c8X[0] - 1;
				lane6c9X[0] <= lane6c9X[0] - 1;
				lane6c10X[0] <= lane6c10X[0] - 1;
				lane6c11X[0] <= lane6c11X[0] - 1;
				lane6c12X[0] <= lane6c12X[0] - 1;
			end
	end
//

/////lane7 control /////
always @(posedge update)
	begin
		if (rst == 1'b1)
			begin //starting position of lane7 cars				
				lane7c0X[0] <= 20;
				lane7c0Y[0] <= 224;
				lane7c1X[0] <= 115;
				lane7c1Y[0] <= 224;
				lane7c2X[0] <= 200;
				lane7c2Y[0] <= 224;
				lane7c3X[0] <= 310;
				lane7c3Y[0] <= 224;
				lane7c4X[0] <= 415;
				lane7c4Y[0] <= 224;
				lane7c5X[0] <= 570;
				lane7c5Y[0] <= 224;
				lane7c6X[0] <= 495;
				lane7c6Y[0] <= 224;
				
			end
			
		//recycling cars back to the start of the lane
		else if (lane7c0X[0] >= 640)
			lane7c0X[0] <= 0;
		else if (lane7c1X[0] >= 640)
			lane7c1X[0] <= 0;
		else if (lane7c2X[0] >= 640)
			lane7c2X[0] <= 0;
		else if (lane7c3X[0] >= 640)
			lane7c3X[0] <= 0;
		else if (lane7c4X[0] >= 640)
			lane7c4X[0] <= 0;
		else if (lane7c5X[0] >= 640)
			lane7c5X[0] <= 0;
		else if (lane7c6X[0] >= 640)
			lane7c6X[0] <= 0;
			
		else
			begin //rate and direction of cars
				lane7c0X[0] <= lane7c0X[0] + 1;
				lane7c1X[0] <= lane7c1X[0] + 1;
				lane7c2X[0] <= lane7c2X[0] + 1;
				lane7c3X[0] <= lane7c3X[0] + 1;
				lane7c4X[0] <= lane7c4X[0] + 1;
				lane7c5X[0] <= lane7c5X[0] + 1;
				lane7c6X[0] <= lane7c6X[0] + 1;
					
			end
	end
//

/////lane8 control /////
always @(posedge update)
	begin
		if (rst == 1'b1)
			begin
				lane8c0X[0] = 300;
				lane8c0Y[0] = 249;
			end
		else if (lane8c0X[0] == 0)
			lane8c0X[0] <= 640;
		else
			lane8c0X[0] <= lane8c0X[0] - 9                                                                                                       ;
	end
//

/////lane9 control /////
always @(posedge update)
	begin
		if (rst == 1'b1)
			begin //starting position of lane9 cars
				lane9c0X[0] <= 30;
				lane9c0Y[0] <= 274;
				lane9c1X[0] <= 150;
				lane9c1Y[0] <= 274;
				lane9c2X[0] <= 255;
				lane9c2Y[0] <= 274;
				lane9c3X[0] <= 365;
				lane9c3Y[0] <= 274;
				lane9c4X[0] <= 465;
				lane9c4Y[0] <= 274;
				lane9c5X[0] <= 570;
				lane9c5Y[0] <= 274;
								
			end
		//recycling cars back to the start of the lane
		else if (lane9c0X[0] >= 640)
			lane9c0X[0] <= 0;
		else if (lane9c1X[0] >= 640)
			lane9c1X[0] <= 0;
		else if (lane9c2X[0] >= 640)
			lane9c2X[0] <= 0;
		else if (lane9c3X[0] >= 640)
			lane9c3X[0] <= 0;
		else if (lane9c4X[0] >= 640)
			lane9c4X[0] <= 0;
		else if (lane9c5X[0] >= 640)
			lane9c5X[0] <= 0;
		
		else
			begin //rate and direction of cars
				lane9c0X[0] <= lane9c0X[0] + 3;
				lane9c1X[0] <= lane9c1X[0] + 3;
				lane9c2X[0] <= lane9c2X[0] + 3;
				lane9c3X[0] <= lane9c3X[0] + 3;
				lane9c4X[0] <= lane9c4X[0] + 3;
				lane9c5X[0] <= lane9c5X[0] + 3;
				
			end
	end
//

/////lane10 control /////
always @(posedge update)
	begin
		if (rst == 1'b1)
			begin //starting position of lane10 cars
				lane10c0X[0] <= 10;
				lane10c0Y[0] <= 299;
				lane10c1X[0] <= 70;
				lane10c1Y[0] <= 299;
				lane10c2X[0] <= 130;
				lane10c2Y[0] <= 299;
				lane10c3X[0] <= 190;
				lane10c3Y[0] <= 299;
				lane10c4X[0] <= 250;
				lane10c4Y[0] <= 299;
				lane10c5X[0] <= 315;
				lane10c5Y[0] <= 299;
				lane10c6X[0] <= 380;
				lane10c6Y[0] <= 299;
				lane10c7X[0] <= 440;
				lane10c7Y[0] <= 299;
				lane10c8X[0] <= 510;
				lane10c8Y[0] <= 299;
				lane10c9X[0] <= 580;
				lane10c9Y[0] <= 299;
								
			end
		//recycling cars back to the start of the lane
		else if (lane10c0X[0] >= 640)
			lane10c0X[0] <= 0;
		else if (lane10c1X[0] >= 640)
			lane10c1X[0] <= 0;
		else if (lane10c2X[0] >= 640)
			lane10c2X[0] <= 0;
		else if (lane10c3X[0] >= 640)
			lane10c3X[0] <= 0;
		else if (lane10c4X[0] >= 640)
			lane10c4X[0] <= 0;
		else if (lane10c5X[0] >= 640)
			lane10c5X[0] <= 0;
		else if (lane10c6X[0] >= 640)
			lane10c6X[0] <= 0;
		else if (lane10c7X[0] >= 640)
			lane10c7X[0] <= 0;
		else if (lane10c8X[0] >= 640)
			lane10c8X[0] <= 0;
		else if (lane10c9X[0] >= 640)
			lane10c9X[0] <= 0;
		
		else
			begin //rate and direction of cars
				lane10c0X[0] <= lane10c0X[0] + 1;
				lane10c1X[0] <= lane10c1X[0] + 1;
				lane10c2X[0] <= lane10c2X[0] + 1;
				lane10c3X[0] <= lane10c3X[0] + 1;
				lane10c4X[0] <= lane10c4X[0] + 1;
				lane10c5X[0] <= lane10c5X[0] + 1;
				lane10c6X[0] <= lane10c6X[0] + 1;
				lane10c7X[0] <= lane10c7X[0] + 1;
				lane10c8X[0] <= lane10c8X[0] + 1;
				lane10c9X[0] <= lane10c9X[0] + 1;
				
			end
	end
//

/////lane11 control /////
always @(posedge update)
	begin
		if (rst == 1'b1)
			begin //starting position of lane11 cars
				lane11c0X[0] <= 30;
				lane11c0Y[0] <= 324;
				lane11c1X[0] <= 100;
				lane11c1Y[0] <= 324;
				lane11c2X[0] <= 170;
				lane11c2Y[0] <= 324;
				lane11c3X[0] <= 240;
				lane11c3Y[0] <= 324;
				lane11c4X[0] <= 310;
				lane11c4Y[0] <= 324;
				lane11c5X[0] <= 385;
				lane11c5Y[0] <= 324;
				lane11c6X[0] <= 450;
				lane11c6Y[0] <= 324;
				lane11c7X[0] <= 520;
				lane11c7Y[0] <= 324;
				lane11c8X[0] <= 580;
				lane11c8Y[0] <= 324;
				
				
			end
		//recycling cars back to the start of the lane
		else if (lane11c0X[0] == 0)
			lane11c0X[0] <= 640;
		else if (lane11c1X[0] == 0)
			lane11c1X[0] <= 640;
		else if (lane11c2X[0] == 0)
			lane11c2X[0] <= 640;
		else if (lane11c3X[0] == 0)
			lane11c3X[0] <= 640;
		else if (lane11c4X[0] == 0)
			lane11c4X[0] <= 640;
		else if (lane11c5X[0] == 0)
			lane11c5X[0] <= 640;
		else if (lane11c6X[0] == 0)
			lane11c6X[0] <= 640;
		else if (lane11c7X[0] == 0)
			lane11c7X[0] <= 640;
		else if (lane11c8X[0] == 0)
			lane11c8X[0] <= 640;
			
		else
			begin //rate and direction of cars
				lane11c0X[0] <= lane11c0X[0] - 1;
				lane11c1X[0] <= lane11c1X[0] - 1;
				lane11c2X[0] <= lane11c2X[0] - 1;
				lane11c3X[0] <= lane11c3X[0] - 1;
				lane11c4X[0] <= lane11c4X[0] - 1;
				lane11c5X[0] <= lane11c5X[0] - 1;
				lane11c6X[0] <= lane11c6X[0] - 1;
				lane11c7X[0] <= lane11c7X[0] - 1;
				lane11c8X[0] <= lane11c8X[0] - 1;
			end
	end
//

/////lane12 control /////
always @(posedge update)
	begin
		if (rst == 1'b1)
			begin //starting position of lane12 cars
				lane12c0X[0] <= 20;
				lane12c0Y[0] <= 349;
				lane12c1X[0] <= 110;
				lane12c1Y[0] <= 349;
				lane12c2X[0] <= 210;
				lane12c2Y[0] <= 349;
				lane12c3X[0] <= 330;
				lane12c3Y[0] <= 349;
				lane12c4X[0] <= 450;
				lane12c4Y[0] <= 349;
				lane12c5X[0] <= 570;
				lane12c5Y[0] <= 349;			
			end
		//recycling cars back to the start of the lane
		else if (lane12c0X[0] == 0)
			lane12c0X[0] <= 640;
		else if (lane12c1X[0] == 0)
			lane12c1X[0] <= 640;
		else if (lane12c2X[0] == 0)
			lane12c2X[0] <= 640;
		else if (lane12c3X[0] == 0)
			lane12c3X[0] <= 640;
		else if (lane12c4X[0] == 0)
			lane12c4X[0] <= 640;
		else if (lane12c5X[0] == 0)
			lane12c5X[0] <= 640;			
		else
			begin //rate and direction of cars
				lane12c0X[0] <= lane12c0X[0] - 2;
				lane12c1X[0] <= lane12c1X[0] - 2;
				lane12c2X[0] <= lane12c2X[0] - 2;
				lane12c3X[0] <= lane12c3X[0] - 2;
				lane12c4X[0] <= lane12c4X[0] - 2;
				lane12c5X[0] <= lane12c5X[0] - 2;
			end
	end
//

/////lane13 control /////
always @(posedge update)
	begin
		if (rst == 1'b1)
			begin //starting position of lane13 cars
				lane13c0X[0] <= 20;
				lane13c0Y[0] <= 374;
				lane13c1X[0] <= 115;
				lane13c1Y[0] <= 374;
				lane13c2X[0] <= 225;
				lane13c2Y[0] <= 374;
				lane13c3X[0] <= 335;
				lane13c3Y[0] <= 374;
				lane13c4X[0] <= 445;
				lane13c4Y[0] <= 374;
				lane13c5X[0] <= 555;
				lane13c5Y[0] <= 374;			
			end
		//recycling cars back to the start of the lane
		else if (lane13c0X[0] >= 640)
			lane13c0X[0] <= 0;
		else if (lane13c1X[0] >= 640)
			lane13c1X[0] <= 0;
		else if (lane13c2X[0] >= 640)
			lane13c2X[0] <= 0;
		else if (lane13c3X[0] >= 640)
			lane13c3X[0] <= 0;
		else if (lane13c4X[0] >= 640)
			lane13c4X[0] <= 0;
		else if (lane13c5X[0] >= 640)
			lane13c5X[0] <= 0;
		else
			begin //rate and direction of cars
				lane13c0X[0] <= lane13c0X[0] + 1;
				lane13c1X[0] <= lane13c1X[0] + 1;
				lane13c2X[0] <= lane13c2X[0] + 1;
				lane13c3X[0] <= lane13c3X[0] + 1;
				lane13c4X[0] <= lane13c4X[0] + 1;
				lane13c5X[0] <= lane13c5X[0] + 1;
			end
	end
//

/////lane14 control /////
always @(posedge update)
	begin
		if (rst == 1'b1)
			begin //starting position of lane14 cars
				lane14c0X[0] <= 24;
				lane14c0Y[0] <= 399;
				lane14c1X[0] <= 150;
				lane14c1Y[0] <= 399;
				lane14c2X[0] <= 290;
				lane14c2Y[0] <= 399;
				lane14c3X[0] <= 440;
				lane14c3Y[0] <= 399;
				lane14c4X[0] <= 570;
				lane14c4Y[0] <= 399;
				
				
			end
		//recycling cars back to the start of the lane
		else if (lane14c0X[0] == 0)
			lane14c0X[0] <= 640;
		else if (lane14c1X[0] == 0)
			lane14c1X[0] <= 640;
		else if (lane14c2X[0] == 0)
			lane14c2X[0] <= 640;
		else if (lane14c3X[0] == 0)
			lane14c3X[0] <= 640;
		else if (lane14c4X[0] == 0)
			lane14c4X[0] <= 640;
			
		else
			begin //rate and direction of cars
				lane14c0X[0] <= lane14c0X[0] - 2;
				lane14c1X[0] <= lane14c1X[0] - 2;
				lane14c2X[0] <= lane14c2X[0] - 2;
				lane14c3X[0] <= lane14c3X[0] - 2;
				lane14c4X[0] <= lane14c4X[0] - 2;
			end
	end
//

/////lane15 control /////
always @(posedge update)
	begin
		if (rst == 1'b1)
			begin //starting position of lane15 cars
				lane15c0X[0] <= 20;
				lane15c0Y[0] <= 424;
				lane15c1X[0] <= 115;
				lane15c1Y[0] <= 424;
				lane15c2X[0] <= 200;
				lane15c2Y[0] <= 424;
				lane15c3X[0] <= 310;
				lane15c3Y[0] <= 424;
				lane15c4X[0] <= 415;
				lane15c4Y[0] <= 424;
				lane15c5X[0] <= 570;
				lane15c5Y[0] <= 424;
				lane15c6X[0] <= 495;
				lane15c6Y[0] <= 424;
				
			end
		//recycling cars back to the start of the lane
		else if (lane15c0X[0] == 0)
			lane15c0X[0] <= 640;
		else if (lane15c1X[0] == 0)
			lane15c1X[0] <= 640;
		else if (lane15c2X[0] == 0)
			lane15c2X[0] <= 640;
		else if (lane15c3X[0] == 0)
			lane15c3X[0] <= 640;
		else if (lane15c4X[0] == 0)
			lane15c4X[0] <= 640;
		else if (lane15c5X[0] == 0)
			lane15c5X[0] <= 640;
		else if (lane15c6X[0] == 0)
			lane15c6X[0] <= 640;
			
		else
			begin //rate and direction of cars
				lane15c0X[0] <= lane15c0X[0] - 1;
				lane15c1X[0] <= lane15c1X[0] - 1;
				lane15c2X[0] <= lane15c2X[0] - 1;
				lane15c3X[0] <= lane15c3X[0] - 1;
				lane15c4X[0] <= lane15c4X[0] - 1;
				lane15c5X[0] <= lane15c5X[0] - 1;
				lane15c6X[0] <= lane15c6X[0] - 1;
			end
	end
//


endmodule 