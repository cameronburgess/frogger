module frogger (board_clk, rst, VGA_R, VGA_G, VGA_B, hsync, vsync, clk, blank_n, up, down, left, right, levelselect);

input board_clk, rst; //, key_clk, keydata; (data from keyboard) 
input up,down,left,right;  //direction inputs from push buttons (3->0 respectively)
input levelselect; //switch that determines the current level
output hsync, vsync, clk, blank_n; //non-color outputs to VGA (including the vga clock "clk", which is the main clock used in this project)

//clocks
clock_converter clocks(board_clk,update,clk); //converts the board clock to VGA clock and frog position update clock (50MHz to 25MHz)
wire clk; //clock that goes to the VGA (primary clock that is used)
wire update; //clock that controls how fast the frog's location updates
//

//frog (player) generator
player_frog	froggy (clk,rst,up,down,left,right,update,xCount,yCount,frog);
wire frog;
//

//car (obstacle) generator
lv1car_generator cars1(clk,update,rst,xCount,yCount,traffic1);
lv2car_generator cars2(clk,update,rst,xCount,yCount,traffic2);
wire [114:0]traffic1;
wire [114:0]traffic2;
//

//level selection
reg [114:0]traffic;

always @(posedge clk)
	begin
		if (levelselect == 1'b0)
			traffic <= traffic1;
		else
			traffic <= traffic2;
	end
//
	
//collision (win/lose condition) calculator	(deal with later)
collision WL(clk,rst,frog,traffic,border,end_zone,xCount,yCount,win,game_over);
wire game_over;
wire win;

//"end zone" that triggers a win - generator
reg end_zone;

always @(posedge clk)
	begin
		end_zone <= ((yCount >= 15) && (yCount <= 65)) ;
	end
//
	
//game area border generator
reg  border;

always @(posedge clk) 
	begin
		border <= (((xCount >= 0) && (xCount < 15) || (xCount >= 630) && (xCount < 641)) || ((yCount >= 0) && (yCount < 15) || (yCount >= 465) && (yCount < 481)));
	end
//

//road line "grid" generator
reg yellow_roadlines;  //between traffic lanes going opposite ways (solid yellow)
reg white_roadlines; //between traffic lanes going the same way (dashed white)

always @(posedge clk)
	begin
		yellow_roadlines <= ( ((yCount >= 69) && (yCount <= 70 )) || ((yCount >= 119) && (yCount <= 120 )) || ((yCount >= 144) && (yCount <= 145 )) || ((yCount >= 169) && (yCount <= 170 )) || ((yCount >= 219) && (yCount <= 220 )) || ((yCount >= 244) && (yCount <= 245 )) || ((yCount >= 269) && (yCount <= 270)) || ((yCount >= 319) && (yCount <= 320 )) || ((yCount >= 369) && (yCount <= 370 )) || ((yCount >= 394) && (yCount <= 395 )) || ((yCount >= 444) && (yCount <= 445 )) );                                                                                                                                                                                                                                                                                                           
		white_roadlines <= (( ((xCount > 15) && (xCount <= 30)) || ((xCount >= 45) && (xCount <= 60)) || ((xCount >= 75) && (xCount <= 90)) || ((xCount >= 105) && (xCount <= 120)) || ((xCount >= 135) && (xCount <= 150)) || ((xCount >= 165) && (xCount <= 180)) || ((xCount >= 195) && (xCount <= 210)) || ((xCount >= 225) && (xCount <= 240)) || ((xCount >= 255) && (xCount <= 270)) || ((xCount >= 285) && (xCount <= 300)) || ((xCount >= 315) && (xCount <= 330)) || ((xCount >= 345) && (xCount <= 360)) || ((xCount >= 375) && (xCount <= 390)) || ((xCount >= 405) && (xCount <= 420)) || ((xCount >= 435) && (xCount <= 450)) || ((xCount >= 465) && (xCount <= 480)) || ((xCount >= 495) && (xCount <= 510)) || ((xCount >= 525) && (xCount <= 540)) || ((xCount >= 555) && (xCount <= 570)) || ((xCount >= 585) && (xCount <= 600)) || ((xCount >= 615) && (xCount < 630)) ) && (((yCount >= 94) && (yCount <= 95 )) || ((yCount >= 194) && (yCount <= 195 )) || ((yCount >= 294) && (yCount <= 295 )) || ((yCount >= 344) && (yCount <= 345 )) || ((yCount >= 419) && (yCount <= 420 )) ));
	end
//

//text/word generator
wire game_over_text;
wire win_text;
wire level_text;
wire level_num1_text;
wire level_num2_text;
wire safezone_L4;
wire safezone_L8;
wire safezone_L13;

text words(clk,rst,xCount,yCount,game_over_text,win_text,level_text,level_num1_text,level_num2_text,safezone_L4,safezone_L8,safezone_L13);
//

//display control
wire [9:0] xCount; 
wire [9:0] yCount;
wire ScreenArea;

VGA_Controller VGA(clk, xCount, yCount, ScreenArea, hsync, vsync, blank_n);

output reg [7:0]VGA_R, VGA_G, VGA_B;

reg R;
reg G;
reg B;

always @(posedge clk)
	begin
		if (game_over == 1'b0)
			begin
				if (win == 1'b0)
					begin;
						if (levelselect == 1'b0)
							begin
								R = (( (border && !level_text && !level_num1_text) || (!frog && safezone_L4) || (!frog && safezone_L8) || (!frog && safezone_L13) || (yellow_roadlines && !frog) || (white_roadlines && !frog) || traffic[0] || traffic [1] || traffic[3] || traffic[4] || traffic[5] || traffic[8] || traffic[9] || traffic[10] || traffic [11] || traffic[13] || traffic[15] || traffic[16] || traffic[17] || traffic[19] || traffic[21] || traffic[22] || traffic[23] || traffic[27] || traffic[28] || traffic[29] || traffic[30] || traffic[32] || traffic[33] || traffic[34] || traffic[35] || traffic[36] || traffic[38] || traffic[40] || traffic[41] || traffic[44] || traffic[45] || traffic[47] || traffic[48] || traffic[50] || traffic[51] || traffic[55] || traffic [56] || traffic[59] || traffic[60] || traffic[62] || traffic[64] || traffic[65] || traffic[67] || traffic[69] || traffic[70] || traffic[72] || traffic[74] || traffic[75] || traffic[77] || traffic[80] || traffic[82] || traffic[84] || traffic[85] || traffic[87] || traffic[89] || traffic[91] || traffic[92] || traffic[94] || traffic[97] || traffic[99] || traffic[101] || traffic[104] || traffic[105] || traffic[106] || traffic[109] || traffic[112] || traffic[113] || traffic[114]));
								G = ((border && !level_text && !level_num1_text) || frog || end_zone || safezone_L4 || safezone_L8 || safezone_L13 || yellow_roadlines || white_roadlines || traffic[9] || traffic[4] || traffic[5] || traffic[6] || traffic[7] || traffic[12] || traffic[13] || traffic[16] || traffic[17] || traffic[18] || traffic[19] || traffic[20] || traffic[21] || traffic[22] || traffic[24] || traffic[25] || traffic[31] || traffic[34] || traffic[35] || traffic[37] || traffic[38] || traffic[40] || traffic[41] || traffic[42] || traffic[44] || traffic[46] || traffic[48] || traffic[49] || traffic[51] || traffic[53] || traffic[55] || traffic[57] || traffic[59] || traffic[61] || traffic[62] || traffic[63] || traffic[65] || traffic[66] || traffic[68] || traffic[70] || traffic[72] || traffic[76] || traffic[77] || traffic[79] || traffic[81] || traffic[82] || traffic[83] || traffic[85] || traffic[86] || traffic[90] || traffic[92] || traffic[93] || traffic[94] || traffic[96] || traffic[98] || traffic[99] || traffic[101] || traffic[102] || traffic[106] || traffic[107] || traffic[108] || traffic[109] || traffic[110] || traffic[113]);
								B = (!frog &&((border && !level_text && !level_num1_text) || end_zone || safezone_L4 || safezone_L8 || safezone_L13 || (white_roadlines && !frog) || traffic[0] || traffic[2] || traffic[3] || traffic[5] || traffic[7] || traffic[11] || traffic[14] || traffic[16] || traffic[20] || traffic[21] || traffic[24] || traffic[26] || traffic[28] || traffic[30] || traffic[31] || traffic[32] || traffic[35] || traffic[39] || traffic[40] || traffic[42] || traffic[43] || traffic[44] || traffic[45] || traffic[46] || traffic[48] || traffic[50] || traffic[52] || traffic[54] || traffic[55] || traffic[57] || traffic[58] || traffic[60] || traffic[61] || traffic[62] || traffic[65] || traffic[67] || traffic[68] || traffic[70] || traffic[71] || traffic[73] || traffic[75] || traffic[77] || traffic[78] || traffic[79] || traffic[82] || traffic[84] || traffic[86] || traffic[88] || traffic[89] || traffic[90] || traffic[91] || traffic[92] || traffic[95] || traffic[96] || traffic[98] || traffic[100] || traffic[101] || traffic[103] || traffic[105] || traffic[107] || traffic[108] || traffic[109] || traffic[111] || traffic[114]));
							end
						else
							begin
								R = (( (border && !level_text && !level_num2_text) || (yellow_roadlines && !frog) || (white_roadlines && !frog) || traffic[0] || traffic [1] || traffic[3] || traffic[4] || traffic[5] || traffic[8] || traffic[9] || traffic[10] || traffic [11] || traffic[13] || traffic[15] || traffic[16] || traffic[17] || traffic[19] || traffic[21] || traffic[22] || traffic[23] || traffic[27] || traffic[28] || traffic[29] || traffic[30] || traffic[32] || traffic[33] || traffic[34] || traffic[35] || traffic[36] || traffic[38] || traffic[40] || traffic[41] || traffic[44] || traffic[45] || traffic[47] || traffic[48] || traffic[50] || traffic[51] || traffic[55] || traffic [56] || traffic[59] || traffic[60] || traffic[62] || traffic[64] || traffic[65] || traffic[67] || traffic[69] || traffic[70] || traffic[72] || traffic[74] || traffic[75] || traffic[77] || traffic[80] || traffic[82] || traffic[84] || traffic[85] || traffic[87] || traffic[89] || traffic[91] || traffic[92] || traffic[94] || traffic[97] || traffic[99] || traffic[101] || traffic[104] || traffic[105] || traffic[106] || traffic[109] || traffic[112] || traffic[113] || traffic[114]));
								G = ((border && !level_text && !level_num2_text) || frog || end_zone || yellow_roadlines || white_roadlines || traffic[9] || traffic[4] || traffic[5] || traffic[6] || traffic[7] || traffic[12] || traffic[13] || traffic[16] || traffic[17] || traffic[18] || traffic[19] || traffic[20] || traffic[21] || traffic[22] || traffic[24] || traffic[25] || traffic[31] || traffic[34] || traffic[35] || traffic[37] || traffic[38] || traffic[40] || traffic[41] || traffic[42] || traffic[44] || traffic[46] || traffic[48] || traffic[49] || traffic[51] || traffic[53] || traffic[55] || traffic[57] || traffic[59] || traffic[61] || traffic[62] || traffic[63] || traffic[65] || traffic[66] || traffic[68] || traffic[70] || traffic[72] || traffic[76] || traffic[77] || traffic[79] || traffic[81] || traffic[82] || traffic[83] || traffic[85] || traffic[86] || traffic[90] || traffic[92] || traffic[93] || traffic[94] || traffic[96] || traffic[98] || traffic[99] || traffic[101] || traffic[102] || traffic[106] || traffic[107] || traffic[108] || traffic[109] || traffic[110] || traffic[113]);
								B = (!frog &&((border && !level_text && !level_num2_text) || end_zone || (white_roadlines && !frog) || traffic[0] || traffic[2] || traffic[3] || traffic[5] || traffic[7] || traffic[11] || traffic[14] || traffic[16] || traffic[20] || traffic[21] || traffic[24] || traffic[26] || traffic[28] || traffic[30] || traffic[31] || traffic[32] || traffic[35] || traffic[39] || traffic[40] || traffic[42] || traffic[43] || traffic[44] || traffic[45] || traffic[46] || traffic[48] || traffic[50] || traffic[52] || traffic[54] || traffic[55] || traffic[57] || traffic[58] || traffic[60] || traffic[61] || traffic[62] || traffic[65] || traffic[67] || traffic[68] || traffic[70] || traffic[71] || traffic[73] || traffic[75] || traffic[77] || traffic[78] || traffic[79] || traffic[82] || traffic[84] || traffic[86] || traffic[88] || traffic[89] || traffic[90] || traffic[91] || traffic[92] || traffic[95] || traffic[96] || traffic[98] || traffic[100] || traffic[101] || traffic[103] || traffic[105] || traffic[107] || traffic[108] || traffic[109] || traffic[111] || traffic[114]));
							end
					end
				else
					begin
						R = 1'b0;
						G = ScreenArea & !win_text;
						B = 1'b0;
					end
			end
		else
			begin
				R = ScreenArea & !game_over_text;
				G = 1'b0;
				B = 1'b0;
			end
	end
//

always@(posedge clk)
	begin
		VGA_R = {8{R}};
		VGA_G = {8{G}};
		VGA_B = {8{B}};
	end 
//

endmodule
